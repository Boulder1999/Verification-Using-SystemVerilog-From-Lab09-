//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
CIM2kEFxO2cMhIAwggn7SyQXXLLSCy+HZj8WVmVRXD3yb2IJ8V8+NgW+XPXIaey/
fYzwDA3KAu7wxaYTLjDtL/d9iHdyiCED2W/ARwziHQz1W4gJXzAJLhOQwrc+4WZE
8WfkSNLkPQTgxJFiXOxm0rWkezbRqKSmAwlKDY3KZK2MHNH9ar+3wDiIBHaJJIsw
1ic4n2txZ0TwZr7XF+P9j5yyB3LbS29I0FG9AmKcTPxzXhubNf0QSz60pnrghAp+
BEWum5szE1gEkPN51tDVuNM7M4i97+TvgHOK6T7TPVHqlV9odrnNY3V9VpfeAOdM
DZ/OU4H6X9clggLaRNa2Bg==
//pragma protect end_key_block
//pragma protect digest_block
svUMM4QUJ/4upu5aMznf0vQhwd4=
//pragma protect end_digest_block
//pragma protect data_block
hqeMKcpFNxcuo2lANSpjNE7/ZKDiVAe2uhSuU95J89YZjvUTSFRGvZ3clnjQSW4W
AYGpJ7vqhLgMLC4+vG37aqlUlbtuTPT9vop9S7lSce+Xfo1YzcNpeUAZNbZ3bsVb
6Mo+yJxOHF6y3JHgbx6+cioSAHqyOLIZFvEYZ+dHpESiU+9Z6FVp0ybr2f3iV32Q
E+3AsUV+9739KFFtxCLo1/aGlD545bVty6wH9ZxKwnmtsQfho0NvsAS/djfF67uJ
4N5psjrk6xZg05FAhqdV1VQvCTd6yI9L28gvXFDF6QdQL28Us9LpW5XIviGP0Jsh
g2c69r1Di/UPWBo3VOLIji8yuMjUDyupCeKRqQkSNryMCKa8D6zZeooOg+d1ltRz
uFZa4quUljavaH4u7Ae/E7KUiAThdp3hBKusOUWbPMpbQJkBqVvPvNWgZeBIfVW3
wWw8e8CYSJs0y7mkZ6uFe47Fc5eGAG28B1oMwAhW31nYiQ19KqKx1WSTpjLSYjPJ
xHTpueELOmQIIYKJGFGa3psjR/sF4Y3XvMnL8Ytu1kPJf3XIoIKAtVOFfaw4MlzS
8zhBkWVl8XGW5tOL2UiX4IFxmWdo4dSH8yI/Fp+C5lwszhzozcmFkFHZpfFgxMLi
6WZ6YUVnQ2M1btgpFuSMYIY6MxnJrLsIILlhPGzNmapDU9CB+ikRevIABnhdDhyP
PqOzK9RPILC4VDpRFZ6D1jdXv1tL00DVlnA480XvpA6d2MC1XOuaCTbUJzijbxJd
hHNXtlgPZndmdbSyoWrBuqWCrGe6NAQ7KXhwoKouBOceM+SycsMGNZDfzuNkN9Lh
aT799hqYVNa4p5FJx8ahV0sKaJ4WxGk2qAOa3jd9BYHcuzj+KpaSgfRxHhfGxHce
b9zO5fyJ5l6WaYoGX9PI7cLQUWhJm2RM7thbAjndpTQMhgtaY7WsOpw+WJtbJ+Bo
Vn3n0o78TUrqgl2sFfYdmteCkmchUZzP5gvCfN1YCzpzGnFnG85TMTAKDHWbh1DV
PRgXb03lhi9duXC/YCscsKXDDNUMO66gHCO5sySr0nvurzGnvdeJhFs9e6VjU4Ei
qwDB7nijfYuVTCLwFYnYULFyMAdvgk28QzJwmslubyJT76Bvv+pMP3auxHT638sm
q7I0wL2aO593B6ucgjO7a2Bqk3/4oUadITp911LDvHjnFxJrxVP4AejffTvUvVq6
+WEIP08TDP8kkCagQNJmL5N/qXdHGO6vmO+Ud9/sLX8uVuP6h/Dp4io2WjNkw7cp
I2aai1YH73xmnMVqGNk1AJCZy66pNDCRQW9g0SJEXPjYxA0xoNQFryzVb4uYTn2y
hrEfhOui2ey2tHB3zYEy/gsmPiXcSL2oO5DK6Mltj1bIi9XBnZvvLJ8lhErtJVPA
2W1KDtPeUnLP7a9GD3tpYL/JjVvOdKImIDil3uSk+C5sy3K92NI99ABF36BQ66J8
i3sW/Q1Wwy0EQPQ+9gvvVRi6Vh0yGnzA3TC9tu32ff9rxvQ8ofiIVB1WxlLUiSOZ
SPfpBIJgSz7r3DaeXt8rQq/ClQhCKEV9uBn/aWAS/SNMkTOTw0Oyy08VNvaPc9pV
Itml232/ruzxq29TpbVEg1GE7wuEfGvoY01OLy8tbe+cfOtqwqvE/mtFv4Edctnh
oIS12vT1LebuC55xlBru3wxuxI2DTzXwaFuB/ncMNbbMvv+swR491pS3CMmL42xr
o7ZkICfE571LxZDUR2pTmd/2Q8muvhcR+egwHsw4vjuV3XdF9veUNsIc7oWZwWo9
2PBwJHR9v4uVe/8DR2E7g/sQGyZ/TphNw7OF43lM97Dv272b2a8a4IfVaIi9vKM+
iFLYxZJvM4ZGbXSiRuu85WoKtqYQ8GHhjjFr/Zsv0TBYA9SLyRaurKT3ASB3tszE
+DdlzB98n69xXy2k4xB8tegVhGzyEJE0NpvfHNDn6fCC9wpYjtuVOl1sStb3nWBt
L33xur2h5sNLEEB70juxuPO2oN7goOgmQ4RQe8YrhcyrgUaixyUFeQ9WD/FRXMTq
zRO8bG/3pOSQEkqh2ilhzBjJ8+KLS+17NjPAYHQ548Dftbxrk3BOgS0ppVrD2AG3
bhQrBJnZrKOyWZWXT2vuRyFE/1cMF2j9sYuuCjRjoxaWk1Bn5M+JA28rRrAB29HY
/nsyjOXk3jnaaEh1HA+6GoCIWwwdqLbdpE+4jYzLQuKCxFnLSRmFJEFpNNunRHOa
FnhVx/eURA7zLS1++O6qB9u9FSOu7sOzuIBvM/g2pVUWiKQ7xpYBoJvQb2pQUsJf
0TSlusRpmoJKBCLYIL/UE+H/D7GNJ3wlTP6gxxGlYcXPFVFjBi2lPj64TubCZ0tY
lEw+cc0lRYCu45m0nD0naPufhZCH1LhI5d6JN3hB73WYwCBbMhCs520Nmp+Xv6N1
HhZ4Js+hGN1djX7xNiwEfVUBnZgD/YGSdpDNaeI54sQAawzwpGAydEehEq6s7Jo1
daCuXpzSbh1VIFKQCibAI55uidD8f8evADRFjfmkzRi2QETDyHcluMvj1EnKvyfk
zSrwjiptTnr+d7YSz3rCphhQZ7qD4RvboNCehmaaj51wSnSX3Oe2HyU9HWXnyG77
3LOdMqi8bf06D+vBbucuihGimxllaJ14L786E0HKqyom5lqBVUFL6I8LOniPFjlC
lAcS31PbBgy5JQiWKQy2tv+/DWcub9ERukezgFONtS5r56WmmmhvDsV4plSGgj05
FRBm/or1X5GxzA8Bq1J1wdFUiUrb8R2KcjeC0+ZUtj/GwFXvJRKeXaF63oKN8r+/
v0i0B9RtXhvJ/cOUnFpCCHcWiuJMlGIpsrKFuY6Wlfky3BAs2649QrvvaUYKvBWN
YY5tTDlDwayK2+nk5l2ZBNh84F/rqldbgpVD7e24Nz0qK49awcVdtmoicxG/EohG
XWOoVAy/yN4191eByoZpXRFco2S5ea1vUaMCZN1K5gZKC2b4Vex6GsNI8whCqkN1
4mN34Qsb1moIWXhSLXNQexX2Bat3nI77/E5vCTq5Oznqm4yiRT2VJkB+LznRZiHP
LlpiGwni7ddyBuPA56J49M4rfmJlbd6af8R5pcEbgrCqIaIF8SNf0fSlmxxMJiLg
VXqJ21paDy8briPzQ5XqRAoIwenkCpoO+T6ljiVJVmAazvFu+YItbhB1/FohGVXZ
6yhUv63XpOqJFgs2oOc3zO8oaNg/NUCW2mFsjiVTypWPcikDy1Pf5G3eoigavsOi
8rLjH8OG3hrBBTZtyKvnLIchfUVRbpC2nDfNK7Xga00QZ+R7gM/2Idf3QybVc5Tq
+PovJiPe5b0QoL0fTyajeO9xnE9TOyb9gkLES/XzPDAhdIyNA7v4fQso8HRquJGn
GKsOG8MzqNKzOc+4nAkWUJ+ZyYQLnR37FQ3zjXnxx2wjBUtG1oY7IxqfSJbQ0zhJ
tQDYifk+Jqp5NduVVjDFh4TEYz7CI9F7l2SSxFhZA2mqUfOHXdLhrNbeBAsVCsDJ
xp0FVA22oKuzrxQDR/mgdAJH8z5alyDfvN3JsPx4O5CDu0AFQFOK2LFEGmmJ7ngc
HZDnpE6EbutYjr6A0oh/OAaqSZ6lU6PXmA1aRFbeI+Mcfgpg1MkNzM9d2UaqmboT
afrXKy3AlZre50K7AFJ206dAzuQzUPDucRmyA83bwF3eaKtgJO1Pi1TjQV22nouV
O8lF3kJb2AOZm+eaWE3g3XVPFMaqyFDRvMtjsAZJy6LLVTwUnCepi33mrakG6mi+
uoEbpdb3w8ShmUmxkv5HnZ6o4/JIic0q/5DCn2TaVA6h0l7IbtOmRwVIs+DrxTAr
S8LZt9aav0wfUyA1ruoiTcYHeh8I3/840Fc/YyO9V/zwW1J1EYz1Oad+jK1HCgxL
AkdV4LTddmiHGMGUx0SW07fYt6iumsGouNukiQJwx8TZmlT85q6tISLj79LlDoUz
60/tthVAY76hYuR+72D/SvKtBtiJz9oHkdCeQafd6fs4gmDgn9BUttvkI86nHQoz
du9B5mgntRRArL7tFlPoih0A5GCjiRmYnpj0Jk1WN7g2UzHePgJUuvbe76DPwKxg
+GgmkSsaFOcHGJmK5OUjt2A/wFf0WFQI5BHcyOGJWxCc6JCtdR0WjZP2rglQ9vk3
VVV2/Cp06+TPOsRw4chK+GfRoaw5vRkIzde6PvjgwCrgRILYeReDrbsqJB+A5FFv
IoI75CRGxraVVHhN00LxBt430eFlr52rVI7BGEvKXB9IaFuqMwCkhbWT4Z54htHV
+xGEyrBEgHGVYKyCfoLfI8gsjGq9EnZsXYuHZwRp8l3EZ5Xv1W4/q99S1jORkjFE
eeJ3gVNSShXkYyTiOZNa+j5KOyEGlWqVCL/qeIMJ5BlPvR5Xi3lxr+EBrDxbauLO
w4NCWL7npArZqS+puQorCSjrua2YqxCShOhRaR5qT6FYDtav9/JscCRg9aPU03Up
2OjSFDlW0ATNiBAiJ4EKw34Gt7tZCjfCW54QPviyEFYglIaRXLWQyV7MLijO+x2y
Bxt6ZI0wMqkFXcVPCcHSOE/jenOUIi+sj2udY+Ev80jjJEXP9XlNQu8Qha0b8ZwI
vvj0i3M7n7gYRqU8Rax0mzO+MU9MjNW++vFjYSfuKuwkFbyHdEns8IPraGnMJbL+
ktLfgwpddplFYUe4bjhqSfXnFvZypeqxUkV2MzXQtdkDUYlwHTAX6/zsrSCmS9sj
wTH/a8csf16b+HRaLGJ+n9QRqXkG6T7qTbgf42Fm0s0IIv5yGMvj0rRahL3VwHYC
2XEcKzyit3waqIm+kVfBP/V3yXbp6UPOrt1WzTk3R63I6zaGeXrX0Ll+S1A5c2WZ
yQlEAprk5ze79c9kGJPYWkTdWKs3RrhbkdKEF1XOr5kFV4Y5LAnOSYdm7jnpywyu
mqQuhYhN91atHa4w2WVKwB31m2ue7nBR8VH6ceOXfXvOFmXe2ktWC+K04bU8m5cp
vz3mVEK+htD/5DvnUVzVCZwYvg3gpCAzvWbQfSwrEHphhd9BLQRirpw3Gb+5ncGY
eSVenW6KoBPYlj9Ws7iF6+5rI7qtuOBvogcJgGZejDhQ7hDJpHAxg2WwTjbU/QqH
QCtXTRf2qs6T9ojXyfS9I/Pb/Bq+odVMbAbJcXKM4vpUlzuLhJA4C2Z3kZbYPIzr
4ni1lw0LY/ARYrNS63rMbyVt1SilzjVctNooHIZa5xxx4fPnL+C3SwcxwL8lXmlT
d3EYW6S5d8ZtohMDqgtp1s8GCAp4VYyCHxQ/Dke1vjaOMxIiE6eY6qtglZhzyVU5
UNs1y/7+/o2zB6AomlKp0kJzJHWegsHhrZdyHI9cGfWSIg8/3niy5owbgvGzG8Eu
RS8VYc8kTPu5gEJ8MbUELco1RqJTWbobL/FyZUX+be2IwaRihZm2if2MnCbiIdL2
cIsLAb11p19eS+0Yk7gyfItkW1cSsIBUf5gIAcWuQsGdZLQF2bCwsCdoHNh3cK7G
ht379JikhBenvQbo554iLT77Y0crTq9RCzIEs+uyY1gro9kyNXHKJiTExD0kZiv3
uR3nnBYN33FAyOBGL5DLZKSZbvJkxNIqxRCLuTDY9MOHHjaKw5YxSjgNACmQL16t
PyJjaxQEYBIFXkYfcZ8ST0AP1oxHthZASIPZEq9IeLIZBFoPT0VDAkY74OCSYP3N
vDdoXqH2fKT8v5ZfgMTuX+/Lx0/tmPVv3gTeR507AjCzM44Dlt1eaG8gquhKwRdJ
UpQmgkA6KmDYoNQdWt71iJLG4q4zfKziVLwwsG1JLMkXsfpke7c6ZEfC3AEYuUaw
r+YK8Px0ynu7wguPUnWOyZbo+NxbTdmBqx/zEN9NDjg1uI69yNtBikJWTtUm61Ah
nlCJx8FAOcTpUSJx88GBzv0DS3fjdI7w8HtDN62/2z+UoNnZbxmd6kZMdzD0miV7
Q0/HxqZ0mQysRPP9vGMHurCS9tJntobo5dCZfEfR67Bb036zOXg7Ljlx6XbDpIDp
ydNRTUfXzPTZRZtwi/hzPheqJN7vZPH+h8KeR4TSS+hGx40R0sZeImgirXqnBNcm
WLgYKH0dtKUzpdQuyUj/yPAUU8SPjeKuz30DrZ6PSWr94lKM83MvIhY/7+19zTHF
X3XLU/D5/pcJRi3O+SvbItWCGjhk1GCLX477VKvk36jJYe2F6THOi7BPa+2G24wB
K6/KAqtA7SEB/3yJVX5mH/WTjE/YPEkkxpCeWtEEq5edaX5MwWZTFRRuwCtQoFcV
A3bMewAGwHUsp2xFoG2YGs27m7PwSBcFjSPNyfUCwbSyFDSwmAx0FqlpCJJK4COq
6ri3BQuoxKcd+frcX2wOuF3FPoRBpUlmF3volABysDa8Zy1hZpg8pUSdfhacClFR
TTxXU3TGtjZJjcjZE82fea6OQRxxxkUJ+ocO17peoE7Pv7+XivTOKyvmmJRTeXXD
e2Uqm//UAofZ9nuiO+ODSl5WTI0EPsycTdOpsJ5la3dKiYPWQuZhyYaQxEzzPuFL
72RFfE6ejFeWbJiuZBjBP848XooT1zvtEOQ0SzvjelG2sbmkX6f8EqhgHpPssvEb
bAXbFQCFZkNGL7hRCPxPQwI6by4bEJFxQgykH+7bZZOFSzTy9BVG8lGxSTtLpfzP
ZjixpLVsszDVgtZZNtVp4OF1GYtN12qwsBRvBENNffm41QvjI8NRBEwINwWpEkFR
EHZhS6fDg+/AgBRqmI2PwzKitOARQ6YP3iboP+C5H6F113xkkfKtWka9oUzv3SK4
2GVlT7fAAnIpVQJVYMQUgSDG/NfKoIDVFfyLEkN+FGOb5in41u3Wh8tYmUM1/LC5
tK2uDh9aJvYQKJVug6EIyxjr+qIIY+AoKdmTjqtc8l6BbSFhNXqQ2OYieNeOy0aV
0BmGd2SF9b4LdB+C2qvjOsMHJjNW8RS1uHDXy6ufNzGAmLznS1myDhREB/buWhKL
ibg4Rzn8IRd74mNpO3y2fj1hqnU77SKeLfQqyOIoJjcY2BNyqDgoiCQSdGkNEhdf
2rGdmeKCsyeirsIyu21+W1Dlx0LVvqludldtGcOosN+85VhWE6wzBSQR0+54tJ/L
MDwRqs5GJMTJ6ikOhsUErjJXHQLeZSgHAMbuE/Wia6Rth1VsUjCt7S6OPrHjajcl
pFplDzUAYB05Vnrv9l8l21163Z8ieLovxuJQAmRjpPCAI1ECqKqJ5qV6MhaTFb9l
bsntE20CYHypitfzHTPfXts/FgUsMRQvL6RkPbveTmYQO0SkcA5kJnntABw2u5zF
RJDJyREL3lTfjKfHcvBLBM9lRxvrVJ+fIeexfyVQGacqG92QiX5vVHJXME9MPVsf
ziL8q/OK5OnnDZtYC6+nHVpePY63pxaeNLdimM2RZU39sLuVBx+sYne5UPrhLWXJ
7Ez4HoG8raW28+NAeZkS3b1IMLTIv4mYLZGNMn9BczFJ+kGXcFg/hWpQF6xp9rZ7
DfF/jSR95LUbDcGRgPdIscvM4X1belqlIjAWnkmo7fzQ4BugDx9LJdQxR+2p7F2Y
G3CE3UXQsBIVG53YeiNO2kGPi/e8ygQFOnFjDgbvHtrxStElFjBJNsxKIpepJI9X
YvjeW+EzsLV8YKoBy/hRWTtsPgiK/lLJNLIvTynX0pJ6fd0JsnPbaoCxFCldVHXV
HF+o89jW8WytQ1BCGmu6ReBd+R4ZcqnJGySAeMHp5OGyhLNhBjZ3Ddp0ztaPbXUR
VRY4nnDhyKbXFAzbRVOMpreUEkdabDzYbYHm4z9NUyGIsp91c1Q1fr1cGsgdRylu
qjUvUOv3ozekjgsjx+NiiKXiJY8kVugIeyTvAL5WCy4cVj2hHkYSOn1uSPp69WBR
TbZTEUiRVItPSBc7CwSUa2R2a0rrxEu1pflTbhVfB0f4V4uEBo5CzymBGcQa8e9p
WsNVl0hTYfQOFSjmmY1XAYwQZ3xWHFP3ndd8zedBkOHttnUHM3n8CrJILt6xJ5JW
k7yaHhFLbNkBdqpn+FO8GZWq8h4+DpvrHkIzhsrmXG5YAnbZmKG7hi2tUNrmOIYu
zXvlJRHWpu1l6WjvjjOzWnvBej0+frppXKFSGACPfhEhRYcc3f45pEhf8mpuWIkg
jaT+qGvGBDPd1zIG18A9psgDNkq7/rW6h6xYDJp3EUiraj9NGijqTQiJfwTzcdw3
uJCNXdc6gjfbSpvxg2nmIRTyfvkckXzBJNG7/6O0Mz5rpl5sBJ8SoKbnRN035Wjo
2M6ewGvLoW7pQ5BwlzzrCGeKWxLiLE7wceXMeRXPbI+2SnT45c38Vno7ya2WheNV
dn1grYd+UJeJ33POkEYvvA3lIQI+DEXYgaZG7FebpGCnitdykQauayXhrkuXCAVz
mOuxJHIxcpFmcBU47HrlHlP36mDOfDDv+9L30Cm6UJZzIbKgcajvlWUI7NpCoL0f
Na7eWqPz1sFcgbxaThzlugYXN2IWW/3bNmynQDR33GXPPQX2BMqk5fE7NbaE0kXZ
6NrPm+KOeprf9dQ9kXJiRbcJjbIfJhOHrqSyEN/S0yhLorTjPbzhDmNm+ju84h6T
OssL7UIxj0cgOuK50tgrIqJY18y5z79SYEQyHRsqjA+C5/g46FWZu23zOjZpYPWx
l5YPlISoDv3o7sxmLKofaf2wMNSxJ4jKq1tnF4VpnOksHuwsJ2IBN4ss8MBy7qfK
wdGEE0hpviYg0YDs3UAiLTRWgRWlJVcRq0m1BCv6QKDI9359BG/CfDPO2EP/l6UY
qpjG/CqWkGjWcgVBudEd/GPQinS7zpDDJywqeFqD+hp/HX0UKxVZgmN5UwVsym6T
XzfmNcPf76LOUR0yFq8VjbLF8Bdp1nY5+wFB3RB4DMPXI+HAaXWGPu1Kwge1LmiB
uRRiFUrCwSK3xGNHiQQYDiFKGCy/Jf1rZtyrqAJPiWcVMACGfmvpwYKRd0UsTCgQ
r9t+bKWnO/gy7nUFe5OPBoJZ0JvoLoTDPBzkYnc3fQkCJ9LDW8X1YpwbUfFyR0xb
CNjE0BoKJJyhRNk7AJxSzZIQmW94yNyG5DTTuM8d18EMS4uKYf88+5NC+DxEn04K
2yRAP/UXJsEiefPpV3D35IjJzQFhVfl4ywGBbUzihWO53BbbV+n9vP8QitNZGoLa
r6UuF6uE7MK68WmVx45AXJGx/eWTCU6NjVb7CwyLYswdXOB2TC7EkjwK9gnVlkss
wM29o8FArw6b2jNqkhKoZRXPcavmxN1q+XUq7BxPsgTBmKoQGyXmJuFoJSx7r/nU
2KRP3NPCNmB/hBRnpDAvn82FGXqqvzwvGc6xJAWZWBbvhjMceC4xogZAl1IdTq66
5bf7XnFpHGrWg2p6H898sx4oG+fS5n2t+6XbWnERQLSmBpvBDq4NlKCRMMKcyIAl
VqnOt7bZqaCqbX4V2ny2p1TUJPsEfFbKLu0V0p/0DQ6MqGsM+hcz4fPFiy0M7yAr
UGy2iJzkhXkOJNYfmW0S/OMjoYKoY/Ny/3ouyulguTEld4uIom1b7f3UkoYCKSqa
npgZME8cBTl8aMwmeAAh9pgOgSiuvgvHsbrdfg0XK3n6gI4ifzftyEffG/gUStJQ
25+dAgpBQt5mN43LYonpE0p0q52C5SwxhhrmbcRTu6kAaK/Mfpei7KVkJ2aqhP3L
hBghMzkXtXx1eXZh7JqeYXGezD7IxuhPalVTsMEEtCLHkGVgZt9AmHiceuT8dbU5
4HxIxkNDe/7Uuq6mbeNmpfnLJX0aEQ4sq/LMzHZ6ZC4k/HSaX65PxH5ZzwyADlBo
AOXycjo3aEbm3d9f4b8jNKugP2A7idS6fNunG9mivy4uaMpX/ZsjSsxk6edLVijd
WPVJfQH7nDcRhuNpogFYnRqY7DdlQddnF2C5VnC7YV2oiWkvG+fbVmT7QztdegeE
EWBy5SNaBENl/WhoZsfhOIHUfm6ithuzpO4+coTB91lV1p+B0ISXE+fyiiEnPBix
l/qg3K8RealUfHOufrJEDGLf27WARmnCi68FaM0kj45uXOrnqLJI4cPajEOSXq10
jNe/Jw2Tx6MwQWz4567kX8uD8MPEsyZSWj4laH6KsoXy2VdYsHyhInCWSvdMAAUo
IXsdJiJJylAOL5A6PU1faojdBRXhD+vsoui3I8CrrKBe7/rftbsOUNYpKL0uot6/
R1wYMoqZKfM6RXk9IefL27TqqmLfhoQwoo6oPH30wBDAdfndPMlxR7rliXicPTMb
//pragma protect end_data_block
//pragma protect digest_block
vd2uzgXny6v8lRzGYynMSJWW6Zw=
//pragma protect end_digest_block
//pragma protect end_protected
